//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "AluAdvance.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [7:0] b;    //: /sn:0 {0}(622,170)(622,134)(#:428,134){1}
//: {2}(426,132)(426,109)(439,109){3}
//: {4}(443,109)(499,109){5}
//: {6}(503,109)(602,109)(#:602,70){7}
//: {8}(501,107)(501,62){9}
//: {10}(441,107)(441,52){11}
//: {12}(424,134)(218,134)(218,164){13}
reg add_switch;    //: /sn:0 {0}(641,268)(641,306){1}
reg carry_in;    //: /sn:0 {0}(630,184)(668,184){1}
reg mul_switch;    //: /sn:0 {0}(285,275)(285,307){1}
reg [7:0] a;    //: /sn:0 {0}(#:202,66)(202,107)(284,107){1}
//: {2}(288,107)(358,107){3}
//: {4}(362,107)(378,107)(378,142){5}
//: {6}(380,144)(590,144)(590,170){7}
//: {8}(#:376,144)(186,144)(186,164){9}
//: {10}(360,105)(360,54){11}
//: {12}(286,105)(286,62){13}
wire carry_out;    //: /sn:0 {0}(551,166)(551,184)(582,184){1}
wire [7:0] add;    //: /sn:0 {0}(#:497,194)(497,229)(604,229){1}
//: {2}(#:606,227)(#:606,199){3}
//: {4}(#:606,231)(606,262){5}
//: {6}(604,264)(523,264){7}
//: {8}(606,266)(606,311)(633,311){9}
wire [7:0] output0;    //: /sn:0 {0}(#:649,311)(675,311)(675,382)(431,382){1}
//: {2}(429,380)(#:429,312)(#:293,312){3}
//: {4}(427,382)(376,382){5}
//: {6}(372,382)(308,382){7}
//: {8}(374,384)(374,439){9}
wire [7:0] mul;    //: /sn:0 {0}(#:277,312)(202,312)(202,261){1}
//: {2}(202,257)(202,217){3}
//: {4}(#:204,215)(304,215)(304,193){5}
//: {6}(202,213)(#:202,193){7}
//: {8}(200,259)(112,259){9}
//: enddecls

  //: LED g44 (add) @(497,187) /sn:0 /w:[ 0 ] /type:1
  //: LED g4 (mul) @(105,259) /sn:0 /R:1 /w:[ 9 ] /type:3
  //: joint g8 (output0) @(374, 382) /w:[ 5 -1 6 8 ]
  _GGBUFIF8 #(4, 6) g47 (.Z(output0), .I(mul), .E(mul_switch));   //: @(283,312) /sn:0 /w:[ 3 0 1 ]
  //: joint g3 (b) @(441, 109) /w:[ 4 10 3 -1 ]
  //: joint g2 (a) @(360, 107) /w:[ 4 10 3 -1 ]
  //: LED g39 (a) @(286,55) /sn:0 /w:[ 13 ] /type:1
  //: LED g1 (b) @(441,45) /sn:0 /w:[ 11 ] /type:3
  //: SWITCH g51 (mul_switch) @(285,262) /sn:0 /R:3 /w:[ 0 ] /st:1 /dn:1
  //: LED g49 (carry_out) @(551,159) /sn:0 /w:[ 0 ] /type:0
  //: SWITCH g50 (carry_in) @(686,184) /sn:0 /R:2 /w:[ 1 ] /st:0 /dn:1
  //: joint g6 (mul) @(202, 259) /w:[ -1 2 8 1 ]
  _GGMUL8 #(124) g35 (.A(a), .B(b), .P(mul));   //: @(202,180) /sn:0 /w:[ 9 13 7 ]
  //: joint g7 (add) @(606, 264) /w:[ -1 5 6 8 ]
  //: LED g9 (output0) @(374,446) /sn:0 /R:2 /w:[ 9 ] /type:3
  //: DIP g31 (a) @(202,56) /sn:0 /w:[ 0 ] /st:10 /dn:1
  _GGADD8 #(68, 70, 62, 64) g36 (.A(a), .B(b), .S(add), .CI(carry_in), .CO(carry_out));   //: @(606,186) /sn:0 /w:[ 7 0 3 0 1 ]
  //: joint g41 (b) @(501, 109) /w:[ 6 8 5 -1 ]
  //: joint g54 (output0) @(429, 382) /w:[ 1 2 4 -1 ]
  //: joint g45 (mul) @(202, 215) /w:[ 4 6 -1 3 ]
  //: SWITCH g52 (add_switch) @(641,255) /sn:0 /R:3 /w:[ 0 ] /st:1 /dn:1
  //: joint g42 (a) @(286, 107) /w:[ 2 12 1 -1 ]
  //: LED g40 (b) @(501,55) /sn:0 /w:[ 9 ] /type:1
  //: DIP g34 (b) @(602,60) /sn:0 /w:[ 7 ] /st:12 /dn:1
  _GGBUFIF8 #(4, 6) g46 (.Z(output0), .I(add), .E(add_switch));   //: @(639,311) /sn:0 /w:[ 0 9 1 ]
  //: LED g5 (add) @(516,264) /sn:0 /R:1 /w:[ 7 ] /type:3
  //: joint g38 (a) @(378, 144) /w:[ 6 5 8 -1 ]
  //: LED g43 (mul) @(304,186) /sn:0 /w:[ 5 ] /type:1
  //: LED g0 (a) @(360,47) /sn:0 /w:[ 11 ] /type:3
  //: joint g48 (add) @(606, 229) /w:[ -1 2 1 4 ]
  //: joint g37 (b) @(426, 134) /w:[ 1 2 12 -1 ]
  //: LED g53 (output0) @(301,382) /sn:0 /R:1 /w:[ 7 ] /type:1

endmodule
//: /netlistEnd


//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "AluRegister.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
supply0 enable;    //: /sn:0 {0}(312,423)(388,423){1}
//: {2}(390,421)(390,264){3}
//: {4}(390,260)(390,122)(316,122){5}
//: {6}(388,262)(314,262){7}
//: {8}(390,425)(390,472){9}
reg clear;    //: /sn:0 {0}(316,112)(401,112){1}
//: {2}(403,110)(403,90){3}
//: {4}(403,114)(403,250){5}
//: {6}(401,252)(314,252){7}
//: {8}(403,254)(403,413)(312,413){9}
reg mul_switch_;    //: /sn:0 {0}(624,367)(624,407){1}
reg [7:0] constant_load;    //: /sn:0 {0}(#:726,217)(650,217){1}
//: {2}(648,215)(#:648,190){3}
//: {4}(646,217)(613,217){5}
//: {6}(648,219)(648,260){7}
//: {8}(650,262)(727,262)(#:727,302){9}
//: {10}(646,262)(586,262)(586,302){11}
reg add_switch;    //: /sn:0 {0}(796,368)(796,407){1}
reg r3_switch;    //: /sn:0 {0}(206,419)(236,419){1}
reg r2_select;    //: /sn:0 {0}(311,337)(311,303){1}
reg carry_in;    //: /sn:0 {0}(767,316)(806,316){1}
reg r1_select;    //: /sn:0 {0}(314,198)(314,163){1}
reg r3_select;    //: /sn:0 {0}(311,514)(311,477){1}
reg r1_switch;    //: /sn:0 {0}(240,117)(208,117){1}
reg r2_switch;    //: /sn:0 {0}(203,256)(238,256){1}
wire carry_out;    //: /sn:0 {0}(719,316)(685,316){1}
wire [7:0] add;    //: /sn:0 {0}(#:743,331)(743,410){1}
//: {2}(745,412)(788,412){3}
//: {4}(#:741,412)(703,412)(703,384){5}
//: {6}(743,414)(743,453){7}
wire [7:0] r1;    //: /sn:0 {0}(#:277,128)(277,161){1}
//: {2}(275,163)(245,163){3}
//: {4}(243,161)(243,149)(213,149){5}
//: {6}(#:243,165)(243,188)(217,188){7}
//: {8}(#:277,165)(277,203)(306,203){9}
wire [7:0] r3;    //: /sn:0 {0}(#:273,429)(273,478){1}
//: {2}(271,480)(239,480){3}
//: {4}(237,478)(237,459)(#:213,459){5}
//: {6}(#:237,482)(237,501)(217,501){7}
//: {8}(#:273,482)(273,519)(303,519){9}
wire [7:0] output0;    //: /sn:0 {0}(#:804,412)(845,412)(845,545)(682,545){1}
//: {2}(#:680,543)(680,412)(#:632,412){3}
//: {4}(678,545)(600,545){5}
//: {6}(598,543)(598,495){7}
//: {8}(#:596,545)(531,545){9}
//: {10}(529,543)(529,506){11}
//: {12}(527,545)(143,545)(143,361){13}
//: {14}(145,359)(273,359)(273,408){15}
//: {16}(143,357)(143,220){17}
//: {18}(145,218)(275,218)(275,247){19}
//: {20}(#:143,216)(143,78)(277,78)(277,107){21}
wire [7:0] input0;    //: /sn:0 {0}(#:319,519)(427,519)(427,344){1}
//: {2}(427,340)(427,284){3}
//: {4}(429,282)(470,282){5}
//: {6}(474,282)(510,282){7}
//: {8}(514,282)(552,282){9}
//: {10}(#:556,282)(759,282)(759,302){11}
//: {12}(554,284)(554,302){13}
//: {14}(512,280)(#:512,256){15}
//: {16}(472,280)(472,236){17}
//: {18}(427,280)(427,203)(#:322,203){19}
//: {20}(425,342)(#:319,342){21}
wire [7:0] mul;    //: /sn:0 {0}(#:616,412)(572,412){1}
//: {2}(570,410)(#:570,331){3}
//: {4}(#:568,412)(524,412)(524,384){5}
//: {6}(#:570,414)(570,435)(507,435){7}
wire [7:0] r2;    //: /sn:0 {0}(#:275,268)(275,302){1}
//: {2}(273,304)(242,304){3}
//: {4}(240,302)(240,287)(212,287){5}
//: {6}(#:240,306)(240,326)(214,326){7}
//: {8}(275,306)(275,342)(303,342){9}
//: enddecls

  //: joint g75 (output0) @(143, 359) /w:[ 14 16 -1 13 ]
  //: LED g4 (output0) @(529,499) /sn:0 /w:[ 11 ] /type:3
  //: joint g8 (r3) @(237, 480) /w:[ 3 4 -1 6 ]
  //: LED g3 (r3) @(210,501) /sn:0 /R:1 /w:[ 7 ] /type:3
  //: SWITCH g90 (r2_select) @(311,290) /sn:0 /R:3 /w:[ 1 ] /st:0 /dn:1
  //: LED g2 (r2) @(207,326) /sn:0 /R:1 /w:[ 7 ] /type:3
  //: SWITCH g91 (r3_select) @(311,464) /sn:0 /R:3 /w:[ 1 ] /st:0 /dn:1
  _GGBUFIF8 #(4, 6) g92 (.Z(input0), .I(r2), .E(r2_select));   //: @(309,342) /sn:0 /w:[ 21 9 0 ]
  //: joint g74 (output0) @(598, 545) /w:[ 5 6 8 -1 ]
  //: joint g104 (add) @(743, 412) /w:[ 2 1 4 6 ]
  //: SWITCH g77 (r1_switch) @(191,117) /sn:0 /w:[ 1 ] /st:0 /dn:1
  //: LED g86 (r1) @(206,149) /sn:0 /R:1 /w:[ 5 ] /type:1
  //: LED g1 (mul) @(500,435) /sn:0 /R:1 /w:[ 7 ] /type:3
  //: LED g60 (constant_load) @(733,217) /sn:0 /R:3 /w:[ 0 ] /type:1
  //: joint g82 (clear) @(403, 252) /w:[ -1 5 6 8 ]
  //: LED g70 (input0) @(512,249) /sn:0 /w:[ 15 ] /type:1
  _GGBUFIF8 #(4, 6) g94 (.Z(input0), .I(r1), .E(r1_select));   //: @(312,203) /sn:0 /w:[ 19 9 0 ]
  //: joint g103 (mul) @(570, 412) /w:[ 1 2 4 6 ]
  //: SWITCH g65 (mul_switch_) @(624,354) /sn:0 /R:3 /w:[ 0 ] /st:0 /dn:1
  //: LED g10 (add) @(743,460) /sn:0 /R:2 /w:[ 7 ] /type:3
  _GGBUFIF8 #(4, 6) g64 (.Z(output0), .I(add), .E(add_switch));   //: @(794,412) /sn:0 /w:[ 0 3 1 ]
  _GGREG8 #(10, 10, 20) g72 (.Q(r2), .D(output0), .EN(enable), .CLR(clear), .CK(r2_switch));   //: @(275,257) /sn:0 /w:[ 0 19 7 7 1 ]
  //: joint g6 (r1) @(243, 163) /w:[ 3 4 -1 6 ]
  _GGADD8 #(68, 70, 62, 64) g56 (.A(constant_load), .B(input0), .S(add), .CI(carry_in), .CO(carry_out));   //: @(743,318) /sn:0 /w:[ 9 11 0 0 0 ]
  _GGREG8 #(10, 10, 20) g73 (.Q(r3), .D(output0), .EN(enable), .CLR(clear), .CK(r3_switch));   //: @(273,418) /sn:0 /w:[ 0 15 0 9 1 ]
  //: joint g68 (output0) @(680, 545) /w:[ 1 2 4 -1 ]
  //: LED g58 (carry_out) @(678,316) /sn:0 /R:1 /w:[ 1 ] /type:0
  //: joint g7 (r2) @(240, 304) /w:[ 3 4 -1 6 ]
  //: LED g9 (constant_load) @(606,217) /sn:0 /R:1 /w:[ 5 ] /type:3
  _GGREG8 #(10, 10, 20) g71 (.Q(r1), .D(output0), .EN(enable), .CLR(clear), .CK(r1_switch));   //: @(277,117) /sn:0 /w:[ 0 21 5 0 0 ]
  //: LED g102 (add) @(703,377) /sn:0 /w:[ 5 ] /type:1
  //: joint g98 (input0) @(512, 282) /w:[ 8 14 7 -1 ]
  //: DIP g59 (constant_load) @(648,180) /sn:0 /w:[ 3 ] /st:0 /dn:1
  //: joint g85 (enable) @(390, 262) /w:[ -1 4 6 3 ]
  //: LED g67 (output0) @(598,488) /sn:0 /w:[ 7 ] /type:1
  //: LED g87 (r2) @(205,287) /sn:0 /R:1 /w:[ 5 ] /type:1
  //: GROUND g83 (enable) @(390,478) /sn:0 /w:[ 9 ]
  //: joint g99 (input0) @(427, 282) /w:[ 4 18 -1 3 ]
  //: joint g81 (clear) @(403, 112) /w:[ -1 2 1 4 ]
  //: joint g69 (input0) @(554, 282) /w:[ 10 -1 9 12 ]
  //: SWITCH g66 (add_switch) @(796,355) /sn:0 /R:3 /w:[ 0 ] /st:1 /dn:1
  //: joint g12 (input0) @(472, 282) /w:[ 6 16 5 -1 ]
  //: SWITCH g57 (carry_in) @(824,316) /sn:0 /R:2 /w:[ 1 ] /st:0 /dn:1
  //: joint g84 (enable) @(390, 423) /w:[ -1 2 1 8 ]
  //: joint g5 (output0) @(529, 545) /w:[ 9 10 12 -1 ]
  //: LED g11 (input0) @(472,229) /sn:0 /w:[ 17 ] /type:3
  //: joint g96 (r2) @(275, 304) /w:[ -1 1 2 8 ]
  //: joint g61 (constant_load) @(648, 262) /w:[ 8 7 10 -1 ]
  //: SWITCH g79 (r3_switch) @(189,419) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g78 (r2_switch) @(186,257) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g97 (r3) @(273, 480) /w:[ -1 1 2 8 ]
  _GGBUFIF8 #(4, 6) g93 (.Z(input0), .I(r3), .E(r3_select));   //: @(309,519) /sn:0 /w:[ 0 9 0 ]
  //: joint g100 (input0) @(427, 342) /w:[ -1 2 20 1 ]
  _GGBUFIF8 #(4, 6) g63 (.Z(output0), .I(mul), .E(mul_switch_));   //: @(622,412) /sn:0 /w:[ 3 0 1 ]
  //: LED g101 (mul) @(524,377) /sn:0 /w:[ 5 ] /type:1
  //: SWITCH g89 (r1_select) @(314,150) /sn:0 /R:3 /w:[ 1 ] /st:1 /dn:1
  //: LED g0 (r1) @(210,188) /sn:0 /R:1 /w:[ 7 ] /type:3
  //: joint g62 (constant_load) @(648, 217) /w:[ 1 2 4 6 ]
  //: SWITCH g80 (clear) @(403,77) /sn:0 /R:3 /w:[ 3 ] /st:0 /dn:1
  //: joint g95 (r1) @(277, 163) /w:[ -1 1 2 8 ]
  //: LED g88 (r3) @(206,459) /sn:0 /R:1 /w:[ 5 ] /type:1
  _GGMUL8 #(1) g55 (.A(input0), .B(constant_load), .P(mul));   //: @(570,318) /sn:0 /delay:" 1" /w:[ 13 11 3 ]
  //: joint g76 (output0) @(143, 218) /w:[ 18 20 -1 17 ]

endmodule
//: /netlistEnd


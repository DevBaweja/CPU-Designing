//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "4bit.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
supply0 enable;    //: /sn:0 {0}(122,437)(201,437){1}
//: {2}(203,435)(203,258){3}
//: {4}(203,254)(203,112){5}
//: {6}(203,108)(203,-30)(129,-30){7}
//: {8}(201,110)(127,110){9}
//: {10}(201,256)(125,256){11}
//: {12}(203,439)(203,558){13}
reg clear;    //: /sn:0 {0}(127,100)(214,100){1}
//: {2}(216,98)(216,-38){3}
//: {4}(216,-42)(216,-73)(203,-73){5}
//: {6}(214,-40)(129,-40){7}
//: {8}(216,102)(216,244){9}
//: {10}(214,246)(125,246){11}
//: {12}(216,248)(216,427)(122,427){13}
reg [7:0] instruction;    //: /sn:0 {0}(#:536,-66)(536,-131){1}
//: {2}(536,-132)(536,-174){3}
//: {4}(536,-175)(536,-188){5}
//: {6}(536,-189)(536,-211){7}
//: {8}(536,-212)(536,-247){9}
//: {10}(536,-248)(#:536,-269){11}
reg [3:0] w24;    //: /sn:0 {0}(#:1116,-222)(1116,-179){1}
//: {2}(1118,-177)(1159,-177){3}
//: {4}(1116,-175)(1116,-136)(1031,-136)(1031,-131){5}
reg w8;    //: /sn:0 {0}(-118,-132)(-90,-132){1}
reg carry_in;    //: /sn:0 {0}(1332,162)(1311,162){1}
reg w9;    //: /sn:0 {0}(856,-90)(888,-90){1}
wire [7:0] w13;    //: /sn:0 {0}(#:1063,-80)(1028,-80){1}
//: {2}(1026,-82)(#:1026,-125){3}
//: {4}(1026,-78)(1026,-10){5}
wire r2_a;    //: /sn:0 {0}(121,-129)(121,185){1}
wire [1:0] w6;    //: /sn:0 {0}(#:531,-247)(-66,-247)(-66,-174){1}
//: {2}(-64,-172)(-26,-172){3}
//: {4}(-66,-170)(-66,-145){5}
wire r1_a;    //: /sn:0 {0}(109,-129)(109,46){1}
wire r1_b;    //: /sn:0 {0}(244,-129)(244,24){1}
wire [7:0] w7;    //: /sn:0 {0}(#:1166,243)(1224,243)(1224,257){1}
//: {2}(1226,259)(1336,259)(1336,244)(#:1324,244){3}
//: {4}(1224,261)(1224,588)(1028,588){5}
//: {6}(1026,586)(1026,338){7}
//: {8}(1026,334)(#:1026,6){9}
//: {10}(1024,336)(962,336){11}
//: {12}(1024,588)(863,588){13}
//: {14}(861,586)(861,500){15}
//: {16}(859,588)(#:-107,588)(-107,398){17}
//: {18}(-105,396)(83,396)(#:83,422){19}
//: {20}(-107,394)(-107,222){21}
//: {22}(-105,220)(86,220)(#:86,241){23}
//: {24}(-107,218)(-107,68){25}
//: {26}(-105,66)(88,66)(#:88,95){27}
//: {28}(#:-107,64)(-107,-74)(90,-74)(90,-45){29}
wire r3_a;    //: /sn:0 {0}(133,360)(133,-129){1}
wire r3_b;    //: /sn:0 {0}(268,-129)(268,342){1}
wire w4;    //: /sn:0 {0}(918,-74)(918,-59){1}
wire [7:0] input_a;    //: /sn:0 {0}(#:153,531)(369,531)(369,367){1}
//: {2}(369,363)(369,192){3}
//: {4}(369,188)(369,116){5}
//: {6}(371,114)(1091,114){7}
//: {8}(#:1095,114)(1303,114)(1303,148){9}
//: {10}(1093,116)(1093,147){11}
//: {12}(369,112)(369,51)(#:117,51){13}
//: {14}(367,190)(#:129,190){15}
//: {16}(367,365)(#:141,365){17}
wire [1:0] w0;    //: /sn:0 {0}(#:540,-131)(912,-131)(912,-103){1}
wire w3;    //: /sn:0 {0}(906,-74)(906,-17)(1041,-17)(1041,-2)(1031,-2){1}
wire [1:0] decode_input_b;    //: /sn:0 {0}(#:531,-174)(362,-174){1}
//: {2}(358,-174)(262,-174)(262,-158){3}
//: {4}(360,-172)(360,-154){5}
wire [1:0] decode_input_a;    //: /sn:0 {0}(#:531,-188)(183,-188){1}
//: {2}(179,-188)(127,-188)(127,-158){3}
//: {4}(181,-186)(181,-158){5}
wire carry_out;    //: /sn:0 {0}(1263,162)(1239,162){1}
wire [7:0] add;    //: /sn:0 {0}(#:1287,177)(1287,242){1}
//: {2}(1289,244)(1308,244){3}
//: {4}(1287,246)(1287,294){5}
wire [7:0] r4;    //: /sn:0 {0}(#:51,494)(81,494){1}
//: {2}(83,492)(#:83,443){3}
//: {4}(#:83,496)(83,512){5}
//: {6}(85,514)(272,514){7}
//: {8}(83,516)(83,531)(137,531){9}
wire [7:0] r1;    //: /sn:0 {0}(#:56,11)(88,11){1}
//: {2}(90,9)(#:90,-24){3}
//: {4}(#:90,13)(90,27){5}
//: {6}(92,29)(236,29){7}
//: {8}(90,31)(90,51)(101,51){9}
wire [7:0] input_b;    //: /sn:0 {0}(#:1125,147)(1125,90){1}
//: {2}(1127,88)(1271,88)(#:1271,148){3}
//: {4}(1123,88)(398,88){5}
//: {6}(396,86)(396,29)(#:252,29){7}
//: {8}(396,90)(396,167){9}
//: {10}(394,169)(#:264,169){11}
//: {12}(396,171)(396,345){13}
//: {14}(394,347)(#:276,347){15}
//: {16}(396,349)(396,514)(#:288,514){17}
wire [7:0] r3;    //: /sn:0 {0}(#:54,328)(84,328){1}
//: {2}(86,326)(#:86,262){3}
//: {4}(#:86,330)(86,345){5}
//: {6}(88,347)(260,347){7}
//: {8}(86,349)(86,365)(125,365){9}
wire decoding;    //: /sn:0 {0}(665,-6)(622,-6)(622,-234)(89,-234)(89,-216){1}
//: {2}(91,-214)(224,-214)(224,-145)(238,-145){3}
//: {4}(89,-212)(89,-145)(103,-145){5}
wire r3_switch;    //: /sn:0 {0}(-60,-116)(-60,252)(49,252){1}
wire r4_b;    //: /sn:0 {0}(280,509)(280,-129){1}
wire r4_switch;    //: /sn:0 {0}(-48,-116)(-48,433)(46,433){1}
wire r4_a;    //: /sn:0 {0}(145,-129)(145,526){1}
wire w2;    //: /sn:0 {0}(1316,239)(1316,225)(894,225)(894,-6){1}
//: {2}(894,-10)(894,-74){3}
//: {4}(892,-8)(686,-8){5}
wire r1_switch;    //: /sn:0 {0}(53,-35)(-84,-35)(-84,-116){1}
wire r2_switch;    //: /sn:0 {0}(-72,-116)(-72,104)(51,104){1}
wire [3:0] w15;    //: /sn:0 {0}(#:540,-211)(1019,-211){1}
//: {2}(1021,-213)(1021,-264){3}
//: {4}(1021,-209)(1021,-131){5}
wire w5;    //: /sn:0 {0}(1158,238)(1158,194)(930,194)(930,-1){1}
//: {2}(930,-5)(930,-74){3}
//: {4}(928,-3)(686,-3){5}
wire r2_b;    //: /sn:0 {0}(256,-129)(256,164){1}
wire [7:0] mul;    //: /sn:0 {0}(#:1109,176)(1109,241){1}
//: {2}(1111,243)(#:1150,243){3}
//: {4}(1109,245)(1109,278){5}
wire [7:0] r2;    //: /sn:0 {0}(#:52,152)(86,152){1}
//: {2}(88,150)(#:88,116){3}
//: {4}(88,154)(88,167){5}
//: {6}(90,169)(248,169){7}
//: {8}(88,171)(88,190)(113,190){9}
//: enddecls

  _GGDECODER4 #(6, 6) g4 (.I(decode_input_b), .E(decoding), .Z0(r1_b), .Z1(r2_b), .Z2(r3_b), .Z3(r4_b));   //: @(262,-145) /sn:0 /w:[ 3 3 0 0 0 1 ] /ss:0 /do:0
  _GGREG8 #(10, 10, 20) g8 (.Q(r4), .D(w7), .EN(enable), .CLR(clear), .CK(r4_switch));   //: @(83,432) /sn:0 /w:[ 3 19 0 13 1 ]
  assign w0 = instruction[7:6]; //: TAP g44 @(534,-131) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  //: joint g75 (w6) @(-66, -172) /w:[ 2 1 -1 4 ]
  //: DIP g16 (instruction) @(536,-279) /sn:0 /w:[ 11 ] /st:49 /dn:1
  //: LED g3 (r3) @(47,328) /sn:0 /R:1 /w:[ 0 ] /type:3
  //: joint g47 (w7) @(1224, 259) /w:[ 2 1 -1 4 ]
  //: joint g26 (input_a) @(369, 365) /w:[ -1 2 16 1 ]
  _GGBUFIF8 #(4, 6) g17 (.Z(input_b), .I(r3), .E(r3_b));   //: @(266,347) /sn:0 /w:[ 15 7 1 ]
  //: LED g2 (r2) @(45,152) /sn:0 /R:1 /w:[ 0 ] /type:3
  //: joint g30 (r4) @(83, 514) /w:[ 6 5 -1 8 ]
  _GGBUFIF8 #(4, 6) g92 (.Z(input_a), .I(r2), .E(r2_a));   //: @(119,190) /sn:0 /w:[ 15 9 1 ]
  //: joint g23 (w2) @(894, -8) /w:[ -1 2 4 1 ]
  //: LED g74 (w6) @(-19,-172) /sn:0 /R:3 /w:[ 3 ] /type:1
  //: joint g24 (clear) @(216, -40) /w:[ -1 4 6 3 ]
  _GGDECODER4 #(3, 3) g1 (.I(decode_input_a), .E(decoding), .Z0(r1_a), .Z1(r2_a), .Z2(r3_a), .Z3(r4_a));   //: @(127,-145) /sn:0 /delay:" 3 3" /w:[ 3 5 0 0 1 0 ] /ss:0 /do:0
  //: LED g39 (w7) @(861,493) /sn:0 /w:[ 15 ] /type:3
  //: joint g77 (decode_input_b) @(360, -174) /w:[ 1 -1 2 4 ]
  //: joint g29 (r3) @(86, 347) /w:[ 6 5 -1 8 ]
  //: LED g60 (w24) @(1166,-177) /sn:0 /R:3 /w:[ 3 ] /type:1
  //: LED g51 (add) @(1287,301) /sn:0 /R:2 /w:[ 5 ] /type:3
  //: joint g18 (enable) @(203, 437) /w:[ -1 2 1 12 ]
  //: joint g82 (clear) @(216, 100) /w:[ -1 2 1 8 ]
  //: LED g70 (decode_input_a) @(181,-151) /sn:0 /R:2 /w:[ 5 ] /type:1
  //: joint g25 (w7) @(-107, 220) /w:[ 22 24 -1 21 ]
  _GGBUFIF8 #(4, 6) g10 (.Z(input_b), .I(r1), .E(r1_b));   //: @(242,29) /sn:0 /w:[ 7 7 1 ]
  _GGBUFIF8 #(4, 6) g94 (.Z(input_a), .I(r1), .E(r1_a));   //: @(107,51) /sn:0 /w:[ 13 9 1 ]
  //: joint g65 (w13) @(1026, -80) /w:[ 1 2 -1 4 ]
  _GGBUFIF8 #(4, 6) g64 (.Z(w7), .I(add), .E(w2));   //: @(1314,244) /sn:0 /w:[ 3 3 0 ]
  _GGREG8 #(10, 10, 20) g72 (.Q(r2), .D(w7), .EN(enable), .CLR(clear), .CK(r2_switch));   //: @(88,105) /sn:0 /w:[ 3 27 9 0 1 ]
  //: joint g49 (mul) @(1109, 243) /w:[ 2 1 -1 4 ]
  //: LED g6 (r4) @(44,494) /sn:0 /R:1 /w:[ 0 ] /type:3
  //: LED g50 (mul) @(1109,285) /sn:0 /R:2 /w:[ 5 ] /type:3
  assign decode_input_a = instruction[3:2]; //: TAP g7 @(534,-188) /sn:0 /R:2 /w:[ 0 5 6 ] /ss:0
  _GGADD8 #(68, 70, 62, 64) g56 (.A(input_b), .B(input_a), .S(add), .CI(carry_in), .CO(carry_out));   //: @(1287,164) /sn:0 /w:[ 3 9 0 1 0 ]
  _GGREG8 #(10, 10, 20) g73 (.Q(r3), .D(w7), .EN(enable), .CLR(clear), .CK(r3_switch));   //: @(86,251) /sn:0 /w:[ 3 23 11 11 1 ]
  //: LED g58 (carry_out) @(1232,162) /sn:0 /R:1 /w:[ 1 ] /type:0
  //: SWITCH g35 (w8) @(-135,-132) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g9 (w7) @(-107, 396) /w:[ 18 20 -1 17 ]
  //: LED g68 (decode_input_b) @(360,-147) /sn:0 /R:2 /w:[ 5 ] /type:1
  //: joint g31 (r2) @(88, 169) /w:[ 6 5 -1 8 ]
  _GGREG8 #(10, 10, 20) g71 (.Q(r1), .D(w7), .EN(enable), .CLR(clear), .CK(r1_switch));   //: @(90,-35) /sn:0 /w:[ 3 29 7 7 0 ]
  _GGOR2 #(6) g22 (.I0(w5), .I1(w2), .Z(decoding));   //: @(675,-6) /sn:0 /R:2 /w:[ 5 5 0 ]
  //: joint g59 (w7) @(1026, 336) /w:[ -1 8 10 7 ]
  //: joint g85 (enable) @(203, 110) /w:[ -1 6 8 5 ]
  //: LED g67 (w15) @(1021,-271) /sn:0 /w:[ 3 ] /type:1
  //: GROUND g83 (enable) @(203,564) /sn:0 /w:[ 13 ]
  //: joint g99 (input_a) @(369, 114) /w:[ 6 12 -1 5 ]
  assign w13 = {w15, w24}; //: CONCAT g45  @(1026,-126) /sn:0 /R:3 /w:[ 3 5 5 ] /dr:1 /tp:0 /drp:1
  //: LED g41 (instruction) @(536,-59) /sn:0 /R:2 /w:[ 0 ] /type:1
  //: joint g33 (input_b) @(396, 169) /w:[ -1 9 10 12 ]
  //: joint g36 (w5) @(930, -3) /w:[ -1 2 4 1 ]
  //: LED g54 (w7) @(955,336) /sn:0 /R:1 /w:[ 11 ] /type:3
  //: comment g42 @(477,138) /sn:0
  //: /line:""
  //: /line:"Instruction Format"
  //: /line:"opcode"
  //: /line:"add"
  //: /line:"mul "
  //: /line:"1 bit = Most significant bit (7 bit)"
  //: /line:""
  //: /line:"4 registors "
  //: /line:"1 registor requires 2 bit "
  //: /line:"Two registor"
  //: /line:"input a of 2 bit = 3 and 2 bit"
  //: /line:"input b of 2 bit = 1 and 0 bit"
  //: /line:""
  //: /line:"values in registor are given by constant load"
  //: /line:"output is unstored"
  //: /line:""
  //: /line:"add/mul r r r"
  //: /line:"make r anynumber + anynumber"
  //: /end
  //: joint g69 (input_a) @(1093, 114) /w:[ 8 -1 7 10 ]
  assign w15 = instruction[3:0]; //: TAP g40 @(534,-211) /sn:0 /R:2 /w:[ 0 7 8 ] /ss:1
  //: joint g52 (add) @(1287, 244) /w:[ 2 1 -1 4 ]
  //: joint g66 (w15) @(1021, -211) /w:[ -1 2 1 4 ]
  _GGBUFIF8 #(4, 6) g12 (.Z(input_b), .I(r2), .E(r2_b));   //: @(254,169) /sn:0 /w:[ 11 7 1 ]
  //: joint g34 (input_b) @(396, 347) /w:[ -1 13 14 16 ]
  _GGBUFIF8 #(4, 6) g28 (.Z(input_b), .I(r4), .E(r4_b));   //: @(278,514) /sn:0 /w:[ 17 7 0 ]
  //: SWITCH g57 (carry_in) @(1350,162) /sn:0 /R:2 /w:[ 0 ] /st:0 /dn:1
  //: joint g46 (w7) @(1026, 588) /w:[ 5 6 12 -1 ]
  //: joint g5 (input_b) @(1125, 88) /w:[ 2 -1 4 1 ]
  _GGBUFIF8 #(4, 6) g14 (.Z(input_a), .I(r4), .E(r4_a));   //: @(143,531) /sn:0 /w:[ 0 9 1 ]
  //: joint g84 (enable) @(203, 256) /w:[ -1 4 10 3 ]
  //: joint g11 (w7) @(861, 588) /w:[ 13 14 16 -1 ]
  //: joint g96 (r2) @(88, 152) /w:[ -1 2 1 4 ]
  //: joint g19 (clear) @(216, 246) /w:[ -1 9 10 12 ]
  _GGDECODER4 #(1, 1) g21 (.I(w6), .E(w8), .Z0(r1_switch), .Z1(r2_switch), .Z2(r3_switch), .Z3(r4_switch));   //: @(-66,-132) /sn:0 /delay:" 1 1" /w:[ 5 1 1 0 0 0 ] /ss:0 /do:0
  //: joint g61 (w24) @(1116, -177) /w:[ 2 1 -1 4 ]
  //: joint g32 (input_b) @(396, 88) /w:[ 5 6 -1 8 ]
  assign decode_input_b = instruction[1:0]; //: TAP g20 @(534,-174) /sn:0 /R:2 /w:[ 0 3 4 ] /ss:0
  //: joint g78 (decode_input_a) @(181, -188) /w:[ 1 -1 2 4 ]
  //: joint g97 (r3) @(86, 328) /w:[ -1 2 1 4 ]
  _GGBUFIF8 #(4, 6) g93 (.Z(input_a), .I(r3), .E(r3_a));   //: @(131,365) /sn:0 /w:[ 17 9 0 ]
  //: joint g100 (input_a) @(369, 190) /w:[ -1 4 14 3 ]
  _GGBUFIF8 #(4, 6) g63 (.Z(w7), .I(mul), .E(w5));   //: @(1156,243) /sn:0 /w:[ 0 3 0 ]
  //: joint g15 (r4) @(83, 494) /w:[ -1 2 1 4 ]
  //: LED g0 (r1) @(49,11) /sn:0 /R:1 /w:[ 0 ] /type:3
  _GGDECODER4 #(6, 6) g43 (.I(w0), .E(w9), .Z0(w2), .Z1(w3), .Z2(w4), .Z3(w5));   //: @(912,-90) /sn:0 /w:[ 1 1 3 0 0 3 ] /ss:0 /do:0
  _GGBUFIF8 #(4, 6) g38 (.Z(w7), .I(w13), .E(w3));   //: @(1026,-4) /sn:0 /R:3 /w:[ 9 5 1 ]
  //: joint g27 (r1) @(90, 29) /w:[ 6 5 -1 8 ]
  //: DIP g48 (w24) @(1116,-232) /sn:0 /w:[ 0 ] /st:5 /dn:1
  //: joint g37 (decoding) @(89, -214) /w:[ 2 1 -1 4 ]
  //: LED g62 (w13) @(1070,-80) /sn:0 /R:3 /w:[ 0 ] /type:1
  //: SWITCH g80 (clear) @(186,-73) /sn:0 /w:[ 5 ] /st:1 /dn:1
  //: joint g95 (r1) @(90, 11) /w:[ -1 2 1 4 ]
  _GGMUL8 #(124) g55 (.A(input_a), .B(input_b), .P(mul));   //: @(1109,163) /sn:0 /w:[ 11 0 0 ]
  //: joint g76 (w7) @(-107, 66) /w:[ 26 28 -1 25 ]
  assign w6 = instruction[5:4]; //: TAP g13 @(534,-247) /sn:0 /R:2 /w:[ 0 9 10 ] /ss:0
  //: SWITCH g53 (w9) @(839,-90) /sn:0 /w:[ 0 ] /st:1 /dn:1

endmodule
//: /netlistEnd

